module part2(); 

endmodule