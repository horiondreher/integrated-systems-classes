// PLL25Hz.v

// Generated using ACDS version 13.1 182 at 2014.04.30.17:06:30

`timescale 1 ps / 1 ps
module PLL25Hz (
		input  wire  clk_in_clk,      //      clk_in.clk
		input  wire  reset_reset,     //       reset.reset
		output wire  clk_out_25m_clk, // clk_out_25m.clk
		input  wire  areset_export,   //      areset.export
		output wire  clk_menor_clk,   //   clk_menor.clk
		output wire  clk_menor2_clk   //  clk_menor2.clk
	);

	PLL25Hz_altpll_0 altpll_0 (
		.clk       (clk_in_clk),      //       inclk_interface.clk
		.reset     (reset_reset),     // inclk_interface_reset.reset
		.read      (),                //             pll_slave.read
		.write     (),                //                      .write
		.address   (),                //                      .address
		.readdata  (),                //                      .readdata
		.writedata (),                //                      .writedata
		.c0        (clk_out_25m_clk), //                    c0.clk
		.c1        (clk_menor_clk),   //                    c1.clk
		.c2        (clk_menor2_clk),  //                    c2.clk
		.areset    (areset_export),   //        areset_conduit.export
		.locked    (),                //        locked_conduit.export
		.phasedone ()                 //     phasedone_conduit.export
	);

endmodule
